module font_rom(
    input wire clk,
    input wire [10:0] addr,
    output reg [7:0] data
);

    always @(posedge clk) begin
        case (addr)
            11'd   0: data <= 8'h00;
            11'd   1: data <= 8'h1C;
            11'd   2: data <= 8'h22;
            11'd   3: data <= 8'h2A;
            11'd   4: data <= 8'h2E;
            11'd   5: data <= 8'h2C;
            11'd   6: data <= 8'h20;
            11'd   7: data <= 8'h1E;
            11'd   8: data <= 8'h00;
            11'd   9: data <= 8'h08;
            11'd  10: data <= 8'h14;
            11'd  11: data <= 8'h22;
            11'd  12: data <= 8'h22;
            11'd  13: data <= 8'h3E;
            11'd  14: data <= 8'h22;
            11'd  15: data <= 8'h22;
            11'd  16: data <= 8'h00;
            11'd  17: data <= 8'h3C;
            11'd  18: data <= 8'h22;
            11'd  19: data <= 8'h22;
            11'd  20: data <= 8'h3C;
            11'd  21: data <= 8'h22;
            11'd  22: data <= 8'h22;
            11'd  23: data <= 8'h3C;
            11'd  24: data <= 8'h00;
            11'd  25: data <= 8'h1C;
            11'd  26: data <= 8'h22;
            11'd  27: data <= 8'h20;
            11'd  28: data <= 8'h20;
            11'd  29: data <= 8'h20;
            11'd  30: data <= 8'h22;
            11'd  31: data <= 8'h1C;
            11'd  32: data <= 8'h00;
            11'd  33: data <= 8'h3C;
            11'd  34: data <= 8'h22;
            11'd  35: data <= 8'h22;
            11'd  36: data <= 8'h22;
            11'd  37: data <= 8'h22;
            11'd  38: data <= 8'h22;
            11'd  39: data <= 8'h3C;
            11'd  40: data <= 8'h00;
            11'd  41: data <= 8'h3E;
            11'd  42: data <= 8'h20;
            11'd  43: data <= 8'h20;
            11'd  44: data <= 8'h3C;
            11'd  45: data <= 8'h20;
            11'd  46: data <= 8'h20;
            11'd  47: data <= 8'h3E;
            11'd  48: data <= 8'h00;
            11'd  49: data <= 8'h3E;
            11'd  50: data <= 8'h20;
            11'd  51: data <= 8'h20;
            11'd  52: data <= 8'h3C;
            11'd  53: data <= 8'h20;
            11'd  54: data <= 8'h20;
            11'd  55: data <= 8'h20;
            11'd  56: data <= 8'h00;
            11'd  57: data <= 8'h1E;
            11'd  58: data <= 8'h20;
            11'd  59: data <= 8'h20;
            11'd  60: data <= 8'h20;
            11'd  61: data <= 8'h26;
            11'd  62: data <= 8'h22;
            11'd  63: data <= 8'h1E;
            11'd  64: data <= 8'h00;
            11'd  65: data <= 8'h22;
            11'd  66: data <= 8'h22;
            11'd  67: data <= 8'h22;
            11'd  68: data <= 8'h3E;
            11'd  69: data <= 8'h22;
            11'd  70: data <= 8'h22;
            11'd  71: data <= 8'h22;
            11'd  72: data <= 8'h00;
            11'd  73: data <= 8'h1C;
            11'd  74: data <= 8'h08;
            11'd  75: data <= 8'h08;
            11'd  76: data <= 8'h08;
            11'd  77: data <= 8'h08;
            11'd  78: data <= 8'h08;
            11'd  79: data <= 8'h1C;
            11'd  80: data <= 8'h00;
            11'd  81: data <= 8'h02;
            11'd  82: data <= 8'h02;
            11'd  83: data <= 8'h02;
            11'd  84: data <= 8'h02;
            11'd  85: data <= 8'h02;
            11'd  86: data <= 8'h22;
            11'd  87: data <= 8'h1C;
            11'd  88: data <= 8'h00;
            11'd  89: data <= 8'h22;
            11'd  90: data <= 8'h24;
            11'd  91: data <= 8'h28;
            11'd  92: data <= 8'h30;
            11'd  93: data <= 8'h28;
            11'd  94: data <= 8'h24;
            11'd  95: data <= 8'h22;
            11'd  96: data <= 8'h00;
            11'd  97: data <= 8'h20;
            11'd  98: data <= 8'h20;
            11'd  99: data <= 8'h20;
            11'd 100: data <= 8'h20;
            11'd 101: data <= 8'h20;
            11'd 102: data <= 8'h20;
            11'd 103: data <= 8'h3E;
            11'd 104: data <= 8'h00;
            11'd 105: data <= 8'h22;
            11'd 106: data <= 8'h36;
            11'd 107: data <= 8'h2A;
            11'd 108: data <= 8'h2A;
            11'd 109: data <= 8'h22;
            11'd 110: data <= 8'h22;
            11'd 111: data <= 8'h22;
            11'd 112: data <= 8'h00;
            11'd 113: data <= 8'h22;
            11'd 114: data <= 8'h22;
            11'd 115: data <= 8'h32;
            11'd 116: data <= 8'h2A;
            11'd 117: data <= 8'h26;
            11'd 118: data <= 8'h22;
            11'd 119: data <= 8'h22;
            11'd 120: data <= 8'h00;
            11'd 121: data <= 8'h1C;
            11'd 122: data <= 8'h22;
            11'd 123: data <= 8'h22;
            11'd 124: data <= 8'h22;
            11'd 125: data <= 8'h22;
            11'd 126: data <= 8'h22;
            11'd 127: data <= 8'h1C;
            11'd 128: data <= 8'h00;
            11'd 129: data <= 8'h3C;
            11'd 130: data <= 8'h22;
            11'd 131: data <= 8'h22;
            11'd 132: data <= 8'h3C;
            11'd 133: data <= 8'h20;
            11'd 134: data <= 8'h20;
            11'd 135: data <= 8'h20;
            11'd 136: data <= 8'h00;
            11'd 137: data <= 8'h1C;
            11'd 138: data <= 8'h22;
            11'd 139: data <= 8'h22;
            11'd 140: data <= 8'h22;
            11'd 141: data <= 8'h2A;
            11'd 142: data <= 8'h24;
            11'd 143: data <= 8'h1A;
            11'd 144: data <= 8'h00;
            11'd 145: data <= 8'h3C;
            11'd 146: data <= 8'h22;
            11'd 147: data <= 8'h22;
            11'd 148: data <= 8'h3C;
            11'd 149: data <= 8'h28;
            11'd 150: data <= 8'h24;
            11'd 151: data <= 8'h22;
            11'd 152: data <= 8'h00;
            11'd 153: data <= 8'h1C;
            11'd 154: data <= 8'h22;
            11'd 155: data <= 8'h20;
            11'd 156: data <= 8'h1C;
            11'd 157: data <= 8'h02;
            11'd 158: data <= 8'h22;
            11'd 159: data <= 8'h1C;
            11'd 160: data <= 8'h00;
            11'd 161: data <= 8'h3E;
            11'd 162: data <= 8'h08;
            11'd 163: data <= 8'h08;
            11'd 164: data <= 8'h08;
            11'd 165: data <= 8'h08;
            11'd 166: data <= 8'h08;
            11'd 167: data <= 8'h08;
            11'd 168: data <= 8'h00;
            11'd 169: data <= 8'h22;
            11'd 170: data <= 8'h22;
            11'd 171: data <= 8'h22;
            11'd 172: data <= 8'h22;
            11'd 173: data <= 8'h22;
            11'd 174: data <= 8'h22;
            11'd 175: data <= 8'h1C;
            11'd 176: data <= 8'h00;
            11'd 177: data <= 8'h22;
            11'd 178: data <= 8'h22;
            11'd 179: data <= 8'h22;
            11'd 180: data <= 8'h22;
            11'd 181: data <= 8'h22;
            11'd 182: data <= 8'h14;
            11'd 183: data <= 8'h08;
            11'd 184: data <= 8'h00;
            11'd 185: data <= 8'h22;
            11'd 186: data <= 8'h22;
            11'd 187: data <= 8'h22;
            11'd 188: data <= 8'h2A;
            11'd 189: data <= 8'h2A;
            11'd 190: data <= 8'h36;
            11'd 191: data <= 8'h22;
            11'd 192: data <= 8'h00;
            11'd 193: data <= 8'h22;
            11'd 194: data <= 8'h22;
            11'd 195: data <= 8'h14;
            11'd 196: data <= 8'h08;
            11'd 197: data <= 8'h14;
            11'd 198: data <= 8'h22;
            11'd 199: data <= 8'h22;
            11'd 200: data <= 8'h00;
            11'd 201: data <= 8'h22;
            11'd 202: data <= 8'h22;
            11'd 203: data <= 8'h14;
            11'd 204: data <= 8'h08;
            11'd 205: data <= 8'h08;
            11'd 206: data <= 8'h08;
            11'd 207: data <= 8'h08;
            11'd 208: data <= 8'h00;
            11'd 209: data <= 8'h3E;
            11'd 210: data <= 8'h02;
            11'd 211: data <= 8'h04;
            11'd 212: data <= 8'h08;
            11'd 213: data <= 8'h10;
            11'd 214: data <= 8'h20;
            11'd 215: data <= 8'h3E;
            11'd 216: data <= 8'h00;
            11'd 217: data <= 8'h3E;
            11'd 218: data <= 8'h30;
            11'd 219: data <= 8'h30;
            11'd 220: data <= 8'h30;
            11'd 221: data <= 8'h30;
            11'd 222: data <= 8'h30;
            11'd 223: data <= 8'h3E;
            11'd 224: data <= 8'h00;
            11'd 225: data <= 8'h00;
            11'd 226: data <= 8'h20;
            11'd 227: data <= 8'h10;
            11'd 228: data <= 8'h08;
            11'd 229: data <= 8'h04;
            11'd 230: data <= 8'h02;
            11'd 231: data <= 8'h00;
            11'd 232: data <= 8'h00;
            11'd 233: data <= 8'h3E;
            11'd 234: data <= 8'h06;
            11'd 235: data <= 8'h06;
            11'd 236: data <= 8'h06;
            11'd 237: data <= 8'h06;
            11'd 238: data <= 8'h06;
            11'd 239: data <= 8'h3E;
            11'd 240: data <= 8'h00;
            11'd 241: data <= 8'h00;
            11'd 242: data <= 8'h00;
            11'd 243: data <= 8'h08;
            11'd 244: data <= 8'h14;
            11'd 245: data <= 8'h22;
            11'd 246: data <= 8'h00;
            11'd 247: data <= 8'h00;
            11'd 248: data <= 8'h00;
            11'd 249: data <= 8'h00;
            11'd 250: data <= 8'h00;
            11'd 251: data <= 8'h00;
            11'd 252: data <= 8'h00;
            11'd 253: data <= 8'h00;
            11'd 254: data <= 8'h00;
            11'd 255: data <= 8'h3E;
            11'd 256: data <= 8'h00;
            11'd 257: data <= 8'h00;
            11'd 258: data <= 8'h00;
            11'd 259: data <= 8'h00;
            11'd 260: data <= 8'h00;
            11'd 261: data <= 8'h00;
            11'd 262: data <= 8'h00;
            11'd 263: data <= 8'h00;
            11'd 264: data <= 8'h00;
            11'd 265: data <= 8'h08;
            11'd 266: data <= 8'h08;
            11'd 267: data <= 8'h08;
            11'd 268: data <= 8'h08;
            11'd 269: data <= 8'h08;
            11'd 270: data <= 8'h00;
            11'd 271: data <= 8'h08;
            11'd 272: data <= 8'h00;
            11'd 273: data <= 8'h14;
            11'd 274: data <= 8'h14;
            11'd 275: data <= 8'h14;
            11'd 276: data <= 8'h00;
            11'd 277: data <= 8'h00;
            11'd 278: data <= 8'h00;
            11'd 279: data <= 8'h00;
            11'd 280: data <= 8'h00;
            11'd 281: data <= 8'h14;
            11'd 282: data <= 8'h14;
            11'd 283: data <= 8'h3E;
            11'd 284: data <= 8'h14;
            11'd 285: data <= 8'h3E;
            11'd 286: data <= 8'h14;
            11'd 287: data <= 8'h14;
            11'd 288: data <= 8'h00;
            11'd 289: data <= 8'h08;
            11'd 290: data <= 8'h1E;
            11'd 291: data <= 8'h28;
            11'd 292: data <= 8'h1C;
            11'd 293: data <= 8'h0A;
            11'd 294: data <= 8'h3C;
            11'd 295: data <= 8'h08;
            11'd 296: data <= 8'h00;
            11'd 297: data <= 8'h30;
            11'd 298: data <= 8'h32;
            11'd 299: data <= 8'h04;
            11'd 300: data <= 8'h08;
            11'd 301: data <= 8'h10;
            11'd 302: data <= 8'h26;
            11'd 303: data <= 8'h06;
            11'd 304: data <= 8'h00;
            11'd 305: data <= 8'h10;
            11'd 306: data <= 8'h28;
            11'd 307: data <= 8'h28;
            11'd 308: data <= 8'h10;
            11'd 309: data <= 8'h2A;
            11'd 310: data <= 8'h24;
            11'd 311: data <= 8'h1A;
            11'd 312: data <= 8'h00;
            11'd 313: data <= 8'h08;
            11'd 314: data <= 8'h08;
            11'd 315: data <= 8'h08;
            11'd 316: data <= 8'h00;
            11'd 317: data <= 8'h00;
            11'd 318: data <= 8'h00;
            11'd 319: data <= 8'h00;
            11'd 320: data <= 8'h00;
            11'd 321: data <= 8'h08;
            11'd 322: data <= 8'h10;
            11'd 323: data <= 8'h20;
            11'd 324: data <= 8'h20;
            11'd 325: data <= 8'h20;
            11'd 326: data <= 8'h10;
            11'd 327: data <= 8'h08;
            11'd 328: data <= 8'h00;
            11'd 329: data <= 8'h08;
            11'd 330: data <= 8'h04;
            11'd 331: data <= 8'h02;
            11'd 332: data <= 8'h02;
            11'd 333: data <= 8'h02;
            11'd 334: data <= 8'h04;
            11'd 335: data <= 8'h08;
            11'd 336: data <= 8'h00;
            11'd 337: data <= 8'h08;
            11'd 338: data <= 8'h2A;
            11'd 339: data <= 8'h1C;
            11'd 340: data <= 8'h08;
            11'd 341: data <= 8'h1C;
            11'd 342: data <= 8'h2A;
            11'd 343: data <= 8'h08;
            11'd 344: data <= 8'h00;
            11'd 345: data <= 8'h00;
            11'd 346: data <= 8'h08;
            11'd 347: data <= 8'h08;
            11'd 348: data <= 8'h3E;
            11'd 349: data <= 8'h08;
            11'd 350: data <= 8'h08;
            11'd 351: data <= 8'h00;
            11'd 352: data <= 8'h00;
            11'd 353: data <= 8'h00;
            11'd 354: data <= 8'h00;
            11'd 355: data <= 8'h00;
            11'd 356: data <= 8'h00;
            11'd 357: data <= 8'h08;
            11'd 358: data <= 8'h08;
            11'd 359: data <= 8'h10;
            11'd 360: data <= 8'h00;
            11'd 361: data <= 8'h00;
            11'd 362: data <= 8'h00;
            11'd 363: data <= 8'h00;
            11'd 364: data <= 8'h3E;
            11'd 365: data <= 8'h00;
            11'd 366: data <= 8'h00;
            11'd 367: data <= 8'h00;
            11'd 368: data <= 8'h00;
            11'd 369: data <= 8'h00;
            11'd 370: data <= 8'h00;
            11'd 371: data <= 8'h00;
            11'd 372: data <= 8'h00;
            11'd 373: data <= 8'h00;
            11'd 374: data <= 8'h00;
            11'd 375: data <= 8'h08;
            11'd 376: data <= 8'h00;
            11'd 377: data <= 8'h00;
            11'd 378: data <= 8'h02;
            11'd 379: data <= 8'h04;
            11'd 380: data <= 8'h08;
            11'd 381: data <= 8'h10;
            11'd 382: data <= 8'h20;
            11'd 383: data <= 8'h00;
            11'd 384: data <= 8'h00;
            11'd 385: data <= 8'h1C;
            11'd 386: data <= 8'h22;
            11'd 387: data <= 8'h26;
            11'd 388: data <= 8'h2A;
            11'd 389: data <= 8'h32;
            11'd 390: data <= 8'h22;
            11'd 391: data <= 8'h1C;
            11'd 392: data <= 8'h00;
            11'd 393: data <= 8'h08;
            11'd 394: data <= 8'h18;
            11'd 395: data <= 8'h08;
            11'd 396: data <= 8'h08;
            11'd 397: data <= 8'h08;
            11'd 398: data <= 8'h08;
            11'd 399: data <= 8'h1C;
            11'd 400: data <= 8'h00;
            11'd 401: data <= 8'h1C;
            11'd 402: data <= 8'h22;
            11'd 403: data <= 8'h02;
            11'd 404: data <= 8'h0C;
            11'd 405: data <= 8'h10;
            11'd 406: data <= 8'h20;
            11'd 407: data <= 8'h3E;
            11'd 408: data <= 8'h00;
            11'd 409: data <= 8'h3E;
            11'd 410: data <= 8'h02;
            11'd 411: data <= 8'h04;
            11'd 412: data <= 8'h0C;
            11'd 413: data <= 8'h02;
            11'd 414: data <= 8'h22;
            11'd 415: data <= 8'h1C;
            11'd 416: data <= 8'h00;
            11'd 417: data <= 8'h04;
            11'd 418: data <= 8'h0C;
            11'd 419: data <= 8'h14;
            11'd 420: data <= 8'h24;
            11'd 421: data <= 8'h3E;
            11'd 422: data <= 8'h04;
            11'd 423: data <= 8'h04;
            11'd 424: data <= 8'h00;
            11'd 425: data <= 8'h3E;
            11'd 426: data <= 8'h20;
            11'd 427: data <= 8'h3C;
            11'd 428: data <= 8'h02;
            11'd 429: data <= 8'h02;
            11'd 430: data <= 8'h22;
            11'd 431: data <= 8'h1C;
            11'd 432: data <= 8'h00;
            11'd 433: data <= 8'h0E;
            11'd 434: data <= 8'h10;
            11'd 435: data <= 8'h20;
            11'd 436: data <= 8'h3C;
            11'd 437: data <= 8'h22;
            11'd 438: data <= 8'h22;
            11'd 439: data <= 8'h1C;
            11'd 440: data <= 8'h00;
            11'd 441: data <= 8'h3E;
            11'd 442: data <= 8'h02;
            11'd 443: data <= 8'h04;
            11'd 444: data <= 8'h08;
            11'd 445: data <= 8'h10;
            11'd 446: data <= 8'h10;
            11'd 447: data <= 8'h10;
            11'd 448: data <= 8'h00;
            11'd 449: data <= 8'h1C;
            11'd 450: data <= 8'h22;
            11'd 451: data <= 8'h22;
            11'd 452: data <= 8'h1C;
            11'd 453: data <= 8'h22;
            11'd 454: data <= 8'h22;
            11'd 455: data <= 8'h1C;
            11'd 456: data <= 8'h00;
            11'd 457: data <= 8'h1C;
            11'd 458: data <= 8'h22;
            11'd 459: data <= 8'h22;
            11'd 460: data <= 8'h1E;
            11'd 461: data <= 8'h02;
            11'd 462: data <= 8'h04;
            11'd 463: data <= 8'h38;
            11'd 464: data <= 8'h00;
            11'd 465: data <= 8'h00;
            11'd 466: data <= 8'h00;
            11'd 467: data <= 8'h08;
            11'd 468: data <= 8'h00;
            11'd 469: data <= 8'h08;
            11'd 470: data <= 8'h00;
            11'd 471: data <= 8'h00;
            11'd 472: data <= 8'h00;
            11'd 473: data <= 8'h00;
            11'd 474: data <= 8'h00;
            11'd 475: data <= 8'h08;
            11'd 476: data <= 8'h00;
            11'd 477: data <= 8'h08;
            11'd 478: data <= 8'h08;
            11'd 479: data <= 8'h10;
            11'd 480: data <= 8'h00;
            11'd 481: data <= 8'h04;
            11'd 482: data <= 8'h08;
            11'd 483: data <= 8'h10;
            11'd 484: data <= 8'h20;
            11'd 485: data <= 8'h10;
            11'd 486: data <= 8'h08;
            11'd 487: data <= 8'h04;
            11'd 488: data <= 8'h00;
            11'd 489: data <= 8'h00;
            11'd 490: data <= 8'h00;
            11'd 491: data <= 8'h3E;
            11'd 492: data <= 8'h00;
            11'd 493: data <= 8'h3E;
            11'd 494: data <= 8'h00;
            11'd 495: data <= 8'h00;
            11'd 496: data <= 8'h00;
            11'd 497: data <= 8'h10;
            11'd 498: data <= 8'h08;
            11'd 499: data <= 8'h04;
            11'd 500: data <= 8'h02;
            11'd 501: data <= 8'h04;
            11'd 502: data <= 8'h08;
            11'd 503: data <= 8'h10;
            11'd 504: data <= 8'h00;
            11'd 505: data <= 8'h1C;
            11'd 506: data <= 8'h22;
            11'd 507: data <= 8'h04;
            11'd 508: data <= 8'h08;
            11'd 509: data <= 8'h08;
            11'd 510: data <= 8'h00;
            11'd 511: data <= 8'h08;
            11'd 512: data <= 8'h80;
            11'd 513: data <= 8'h9C;
            11'd 514: data <= 8'hA2;
            11'd 515: data <= 8'hAA;
            11'd 516: data <= 8'hAE;
            11'd 517: data <= 8'hAC;
            11'd 518: data <= 8'hA0;
            11'd 519: data <= 8'h9E;
            11'd 520: data <= 8'h80;
            11'd 521: data <= 8'h88;
            11'd 522: data <= 8'h94;
            11'd 523: data <= 8'hA2;
            11'd 524: data <= 8'hA2;
            11'd 525: data <= 8'hBE;
            11'd 526: data <= 8'hA2;
            11'd 527: data <= 8'hA2;
            11'd 528: data <= 8'h80;
            11'd 529: data <= 8'hBC;
            11'd 530: data <= 8'hA2;
            11'd 531: data <= 8'hA2;
            11'd 532: data <= 8'hBC;
            11'd 533: data <= 8'hA2;
            11'd 534: data <= 8'hA2;
            11'd 535: data <= 8'hBC;
            11'd 536: data <= 8'h80;
            11'd 537: data <= 8'h9C;
            11'd 538: data <= 8'hA2;
            11'd 539: data <= 8'hA0;
            11'd 540: data <= 8'hA0;
            11'd 541: data <= 8'hA0;
            11'd 542: data <= 8'hA2;
            11'd 543: data <= 8'h9C;
            11'd 544: data <= 8'h80;
            11'd 545: data <= 8'hBC;
            11'd 546: data <= 8'hA2;
            11'd 547: data <= 8'hA2;
            11'd 548: data <= 8'hA2;
            11'd 549: data <= 8'hA2;
            11'd 550: data <= 8'hA2;
            11'd 551: data <= 8'hBC;
            11'd 552: data <= 8'h80;
            11'd 553: data <= 8'hBE;
            11'd 554: data <= 8'hA0;
            11'd 555: data <= 8'hA0;
            11'd 556: data <= 8'hBC;
            11'd 557: data <= 8'hA0;
            11'd 558: data <= 8'hA0;
            11'd 559: data <= 8'hBE;
            11'd 560: data <= 8'h80;
            11'd 561: data <= 8'hBE;
            11'd 562: data <= 8'hA0;
            11'd 563: data <= 8'hA0;
            11'd 564: data <= 8'hBC;
            11'd 565: data <= 8'hA0;
            11'd 566: data <= 8'hA0;
            11'd 567: data <= 8'hA0;
            11'd 568: data <= 8'h80;
            11'd 569: data <= 8'h9E;
            11'd 570: data <= 8'hA0;
            11'd 571: data <= 8'hA0;
            11'd 572: data <= 8'hA0;
            11'd 573: data <= 8'hA6;
            11'd 574: data <= 8'hA2;
            11'd 575: data <= 8'h9E;
            11'd 576: data <= 8'h80;
            11'd 577: data <= 8'hA2;
            11'd 578: data <= 8'hA2;
            11'd 579: data <= 8'hA2;
            11'd 580: data <= 8'hBE;
            11'd 581: data <= 8'hA2;
            11'd 582: data <= 8'hA2;
            11'd 583: data <= 8'hA2;
            11'd 584: data <= 8'h80;
            11'd 585: data <= 8'h9C;
            11'd 586: data <= 8'h88;
            11'd 587: data <= 8'h88;
            11'd 588: data <= 8'h88;
            11'd 589: data <= 8'h88;
            11'd 590: data <= 8'h88;
            11'd 591: data <= 8'h9C;
            11'd 592: data <= 8'h80;
            11'd 593: data <= 8'h82;
            11'd 594: data <= 8'h82;
            11'd 595: data <= 8'h82;
            11'd 596: data <= 8'h82;
            11'd 597: data <= 8'h82;
            11'd 598: data <= 8'hA2;
            11'd 599: data <= 8'h9C;
            11'd 600: data <= 8'h80;
            11'd 601: data <= 8'hA2;
            11'd 602: data <= 8'hA4;
            11'd 603: data <= 8'hA8;
            11'd 604: data <= 8'hB0;
            11'd 605: data <= 8'hA8;
            11'd 606: data <= 8'hA4;
            11'd 607: data <= 8'hA2;
            11'd 608: data <= 8'h80;
            11'd 609: data <= 8'hA0;
            11'd 610: data <= 8'hA0;
            11'd 611: data <= 8'hA0;
            11'd 612: data <= 8'hA0;
            11'd 613: data <= 8'hA0;
            11'd 614: data <= 8'hA0;
            11'd 615: data <= 8'hBE;
            11'd 616: data <= 8'h80;
            11'd 617: data <= 8'hA2;
            11'd 618: data <= 8'hB6;
            11'd 619: data <= 8'hAA;
            11'd 620: data <= 8'hAA;
            11'd 621: data <= 8'hA2;
            11'd 622: data <= 8'hA2;
            11'd 623: data <= 8'hA2;
            11'd 624: data <= 8'h80;
            11'd 625: data <= 8'hA2;
            11'd 626: data <= 8'hA2;
            11'd 627: data <= 8'hB2;
            11'd 628: data <= 8'hAA;
            11'd 629: data <= 8'hA6;
            11'd 630: data <= 8'hA2;
            11'd 631: data <= 8'hA2;
            11'd 632: data <= 8'h80;
            11'd 633: data <= 8'h9C;
            11'd 634: data <= 8'hA2;
            11'd 635: data <= 8'hA2;
            11'd 636: data <= 8'hA2;
            11'd 637: data <= 8'hA2;
            11'd 638: data <= 8'hA2;
            11'd 639: data <= 8'h9C;
            11'd 640: data <= 8'h80;
            11'd 641: data <= 8'hBC;
            11'd 642: data <= 8'hA2;
            11'd 643: data <= 8'hA2;
            11'd 644: data <= 8'hBC;
            11'd 645: data <= 8'hA0;
            11'd 646: data <= 8'hA0;
            11'd 647: data <= 8'hA0;
            11'd 648: data <= 8'h80;
            11'd 649: data <= 8'h9C;
            11'd 650: data <= 8'hA2;
            11'd 651: data <= 8'hA2;
            11'd 652: data <= 8'hA2;
            11'd 653: data <= 8'hAA;
            11'd 654: data <= 8'hA4;
            11'd 655: data <= 8'h9A;
            11'd 656: data <= 8'h80;
            11'd 657: data <= 8'hBC;
            11'd 658: data <= 8'hA2;
            11'd 659: data <= 8'hA2;
            11'd 660: data <= 8'hBC;
            11'd 661: data <= 8'hA8;
            11'd 662: data <= 8'hA4;
            11'd 663: data <= 8'hA2;
            11'd 664: data <= 8'h80;
            11'd 665: data <= 8'h9C;
            11'd 666: data <= 8'hA2;
            11'd 667: data <= 8'hA0;
            11'd 668: data <= 8'h9C;
            11'd 669: data <= 8'h82;
            11'd 670: data <= 8'hA2;
            11'd 671: data <= 8'h9C;
            11'd 672: data <= 8'h80;
            11'd 673: data <= 8'hBE;
            11'd 674: data <= 8'h88;
            11'd 675: data <= 8'h88;
            11'd 676: data <= 8'h88;
            11'd 677: data <= 8'h88;
            11'd 678: data <= 8'h88;
            11'd 679: data <= 8'h88;
            11'd 680: data <= 8'h80;
            11'd 681: data <= 8'hA2;
            11'd 682: data <= 8'hA2;
            11'd 683: data <= 8'hA2;
            11'd 684: data <= 8'hA2;
            11'd 685: data <= 8'hA2;
            11'd 686: data <= 8'hA2;
            11'd 687: data <= 8'h9C;
            11'd 688: data <= 8'h80;
            11'd 689: data <= 8'hA2;
            11'd 690: data <= 8'hA2;
            11'd 691: data <= 8'hA2;
            11'd 692: data <= 8'hA2;
            11'd 693: data <= 8'hA2;
            11'd 694: data <= 8'h94;
            11'd 695: data <= 8'h88;
            11'd 696: data <= 8'h80;
            11'd 697: data <= 8'hA2;
            11'd 698: data <= 8'hA2;
            11'd 699: data <= 8'hA2;
            11'd 700: data <= 8'hAA;
            11'd 701: data <= 8'hAA;
            11'd 702: data <= 8'hB6;
            11'd 703: data <= 8'hA2;
            11'd 704: data <= 8'h80;
            11'd 705: data <= 8'hA2;
            11'd 706: data <= 8'hA2;
            11'd 707: data <= 8'h94;
            11'd 708: data <= 8'h88;
            11'd 709: data <= 8'h94;
            11'd 710: data <= 8'hA2;
            11'd 711: data <= 8'hA2;
            11'd 712: data <= 8'h80;
            11'd 713: data <= 8'hA2;
            11'd 714: data <= 8'hA2;
            11'd 715: data <= 8'h94;
            11'd 716: data <= 8'h88;
            11'd 717: data <= 8'h88;
            11'd 718: data <= 8'h88;
            11'd 719: data <= 8'h88;
            11'd 720: data <= 8'h80;
            11'd 721: data <= 8'hBE;
            11'd 722: data <= 8'h82;
            11'd 723: data <= 8'h84;
            11'd 724: data <= 8'h88;
            11'd 725: data <= 8'h90;
            11'd 726: data <= 8'hA0;
            11'd 727: data <= 8'hBE;
            11'd 728: data <= 8'h80;
            11'd 729: data <= 8'hBE;
            11'd 730: data <= 8'hB0;
            11'd 731: data <= 8'hB0;
            11'd 732: data <= 8'hB0;
            11'd 733: data <= 8'hB0;
            11'd 734: data <= 8'hB0;
            11'd 735: data <= 8'hBE;
            11'd 736: data <= 8'h80;
            11'd 737: data <= 8'h80;
            11'd 738: data <= 8'hA0;
            11'd 739: data <= 8'h90;
            11'd 740: data <= 8'h88;
            11'd 741: data <= 8'h84;
            11'd 742: data <= 8'h82;
            11'd 743: data <= 8'h80;
            11'd 744: data <= 8'h80;
            11'd 745: data <= 8'hBE;
            11'd 746: data <= 8'h86;
            11'd 747: data <= 8'h86;
            11'd 748: data <= 8'h86;
            11'd 749: data <= 8'h86;
            11'd 750: data <= 8'h86;
            11'd 751: data <= 8'hBE;
            11'd 752: data <= 8'h80;
            11'd 753: data <= 8'h80;
            11'd 754: data <= 8'h80;
            11'd 755: data <= 8'h88;
            11'd 756: data <= 8'h94;
            11'd 757: data <= 8'hA2;
            11'd 758: data <= 8'h80;
            11'd 759: data <= 8'h80;
            11'd 760: data <= 8'h80;
            11'd 761: data <= 8'h80;
            11'd 762: data <= 8'h80;
            11'd 763: data <= 8'h80;
            11'd 764: data <= 8'h80;
            11'd 765: data <= 8'h80;
            11'd 766: data <= 8'h80;
            11'd 767: data <= 8'hBE;
            11'd 768: data <= 8'h80;
            11'd 769: data <= 8'h80;
            11'd 770: data <= 8'h80;
            11'd 771: data <= 8'h80;
            11'd 772: data <= 8'h80;
            11'd 773: data <= 8'h80;
            11'd 774: data <= 8'h80;
            11'd 775: data <= 8'h80;
            11'd 776: data <= 8'h80;
            11'd 777: data <= 8'h88;
            11'd 778: data <= 8'h88;
            11'd 779: data <= 8'h88;
            11'd 780: data <= 8'h88;
            11'd 781: data <= 8'h88;
            11'd 782: data <= 8'h80;
            11'd 783: data <= 8'h88;
            11'd 784: data <= 8'h80;
            11'd 785: data <= 8'h94;
            11'd 786: data <= 8'h94;
            11'd 787: data <= 8'h94;
            11'd 788: data <= 8'h80;
            11'd 789: data <= 8'h80;
            11'd 790: data <= 8'h80;
            11'd 791: data <= 8'h80;
            11'd 792: data <= 8'h80;
            11'd 793: data <= 8'h94;
            11'd 794: data <= 8'h94;
            11'd 795: data <= 8'hBE;
            11'd 796: data <= 8'h94;
            11'd 797: data <= 8'hBE;
            11'd 798: data <= 8'h94;
            11'd 799: data <= 8'h94;
            11'd 800: data <= 8'h80;
            11'd 801: data <= 8'h88;
            11'd 802: data <= 8'h9E;
            11'd 803: data <= 8'hA8;
            11'd 804: data <= 8'h9C;
            11'd 805: data <= 8'h8A;
            11'd 806: data <= 8'hBC;
            11'd 807: data <= 8'h88;
            11'd 808: data <= 8'h80;
            11'd 809: data <= 8'hB0;
            11'd 810: data <= 8'hB2;
            11'd 811: data <= 8'h84;
            11'd 812: data <= 8'h88;
            11'd 813: data <= 8'h90;
            11'd 814: data <= 8'hA6;
            11'd 815: data <= 8'h86;
            11'd 816: data <= 8'h80;
            11'd 817: data <= 8'h90;
            11'd 818: data <= 8'hA8;
            11'd 819: data <= 8'hA8;
            11'd 820: data <= 8'h90;
            11'd 821: data <= 8'hAA;
            11'd 822: data <= 8'hA4;
            11'd 823: data <= 8'h9A;
            11'd 824: data <= 8'h80;
            11'd 825: data <= 8'h88;
            11'd 826: data <= 8'h88;
            11'd 827: data <= 8'h88;
            11'd 828: data <= 8'h80;
            11'd 829: data <= 8'h80;
            11'd 830: data <= 8'h80;
            11'd 831: data <= 8'h80;
            11'd 832: data <= 8'h80;
            11'd 833: data <= 8'h88;
            11'd 834: data <= 8'h90;
            11'd 835: data <= 8'hA0;
            11'd 836: data <= 8'hA0;
            11'd 837: data <= 8'hA0;
            11'd 838: data <= 8'h90;
            11'd 839: data <= 8'h88;
            11'd 840: data <= 8'h80;
            11'd 841: data <= 8'h88;
            11'd 842: data <= 8'h84;
            11'd 843: data <= 8'h82;
            11'd 844: data <= 8'h82;
            11'd 845: data <= 8'h82;
            11'd 846: data <= 8'h84;
            11'd 847: data <= 8'h88;
            11'd 848: data <= 8'h80;
            11'd 849: data <= 8'h88;
            11'd 850: data <= 8'hAA;
            11'd 851: data <= 8'h9C;
            11'd 852: data <= 8'h88;
            11'd 853: data <= 8'h9C;
            11'd 854: data <= 8'hAA;
            11'd 855: data <= 8'h88;
            11'd 856: data <= 8'h80;
            11'd 857: data <= 8'h80;
            11'd 858: data <= 8'h88;
            11'd 859: data <= 8'h88;
            11'd 860: data <= 8'hBE;
            11'd 861: data <= 8'h88;
            11'd 862: data <= 8'h88;
            11'd 863: data <= 8'h80;
            11'd 864: data <= 8'h80;
            11'd 865: data <= 8'h80;
            11'd 866: data <= 8'h80;
            11'd 867: data <= 8'h80;
            11'd 868: data <= 8'h80;
            11'd 869: data <= 8'h88;
            11'd 870: data <= 8'h88;
            11'd 871: data <= 8'h90;
            11'd 872: data <= 8'h80;
            11'd 873: data <= 8'h80;
            11'd 874: data <= 8'h80;
            11'd 875: data <= 8'h80;
            11'd 876: data <= 8'hBE;
            11'd 877: data <= 8'h80;
            11'd 878: data <= 8'h80;
            11'd 879: data <= 8'h80;
            11'd 880: data <= 8'h80;
            11'd 881: data <= 8'h80;
            11'd 882: data <= 8'h80;
            11'd 883: data <= 8'h80;
            11'd 884: data <= 8'h80;
            11'd 885: data <= 8'h80;
            11'd 886: data <= 8'h80;
            11'd 887: data <= 8'h88;
            11'd 888: data <= 8'h80;
            11'd 889: data <= 8'h80;
            11'd 890: data <= 8'h82;
            11'd 891: data <= 8'h84;
            11'd 892: data <= 8'h88;
            11'd 893: data <= 8'h90;
            11'd 894: data <= 8'hA0;
            11'd 895: data <= 8'h80;
            11'd 896: data <= 8'h80;
            11'd 897: data <= 8'h9C;
            11'd 898: data <= 8'hA2;
            11'd 899: data <= 8'hA6;
            11'd 900: data <= 8'hAA;
            11'd 901: data <= 8'hB2;
            11'd 902: data <= 8'hA2;
            11'd 903: data <= 8'h9C;
            11'd 904: data <= 8'h80;
            11'd 905: data <= 8'h88;
            11'd 906: data <= 8'h98;
            11'd 907: data <= 8'h88;
            11'd 908: data <= 8'h88;
            11'd 909: data <= 8'h88;
            11'd 910: data <= 8'h88;
            11'd 911: data <= 8'h9C;
            11'd 912: data <= 8'h80;
            11'd 913: data <= 8'h9C;
            11'd 914: data <= 8'hA2;
            11'd 915: data <= 8'h82;
            11'd 916: data <= 8'h8C;
            11'd 917: data <= 8'h90;
            11'd 918: data <= 8'hA0;
            11'd 919: data <= 8'hBE;
            11'd 920: data <= 8'h80;
            11'd 921: data <= 8'hBE;
            11'd 922: data <= 8'h82;
            11'd 923: data <= 8'h84;
            11'd 924: data <= 8'h8C;
            11'd 925: data <= 8'h82;
            11'd 926: data <= 8'hA2;
            11'd 927: data <= 8'h9C;
            11'd 928: data <= 8'h80;
            11'd 929: data <= 8'h84;
            11'd 930: data <= 8'h8C;
            11'd 931: data <= 8'h94;
            11'd 932: data <= 8'hA4;
            11'd 933: data <= 8'hBE;
            11'd 934: data <= 8'h84;
            11'd 935: data <= 8'h84;
            11'd 936: data <= 8'h80;
            11'd 937: data <= 8'hBE;
            11'd 938: data <= 8'hA0;
            11'd 939: data <= 8'hBC;
            11'd 940: data <= 8'h82;
            11'd 941: data <= 8'h82;
            11'd 942: data <= 8'hA2;
            11'd 943: data <= 8'h9C;
            11'd 944: data <= 8'h80;
            11'd 945: data <= 8'h8E;
            11'd 946: data <= 8'h90;
            11'd 947: data <= 8'hA0;
            11'd 948: data <= 8'hBC;
            11'd 949: data <= 8'hA2;
            11'd 950: data <= 8'hA2;
            11'd 951: data <= 8'h9C;
            11'd 952: data <= 8'h80;
            11'd 953: data <= 8'hBE;
            11'd 954: data <= 8'h82;
            11'd 955: data <= 8'h84;
            11'd 956: data <= 8'h88;
            11'd 957: data <= 8'h90;
            11'd 958: data <= 8'h90;
            11'd 959: data <= 8'h90;
            11'd 960: data <= 8'h80;
            11'd 961: data <= 8'h9C;
            11'd 962: data <= 8'hA2;
            11'd 963: data <= 8'hA2;
            11'd 964: data <= 8'h9C;
            11'd 965: data <= 8'hA2;
            11'd 966: data <= 8'hA2;
            11'd 967: data <= 8'h9C;
            11'd 968: data <= 8'h80;
            11'd 969: data <= 8'h9C;
            11'd 970: data <= 8'hA2;
            11'd 971: data <= 8'hA2;
            11'd 972: data <= 8'h9E;
            11'd 973: data <= 8'h82;
            11'd 974: data <= 8'h84;
            11'd 975: data <= 8'hB8;
            11'd 976: data <= 8'h80;
            11'd 977: data <= 8'h80;
            11'd 978: data <= 8'h80;
            11'd 979: data <= 8'h88;
            11'd 980: data <= 8'h80;
            11'd 981: data <= 8'h88;
            11'd 982: data <= 8'h80;
            11'd 983: data <= 8'h80;
            11'd 984: data <= 8'h80;
            11'd 985: data <= 8'h80;
            11'd 986: data <= 8'h80;
            11'd 987: data <= 8'h88;
            11'd 988: data <= 8'h80;
            11'd 989: data <= 8'h88;
            11'd 990: data <= 8'h88;
            11'd 991: data <= 8'h90;
            11'd 992: data <= 8'h80;
            11'd 993: data <= 8'h84;
            11'd 994: data <= 8'h88;
            11'd 995: data <= 8'h90;
            11'd 996: data <= 8'hA0;
            11'd 997: data <= 8'h90;
            11'd 998: data <= 8'h88;
            11'd 999: data <= 8'h84;
            11'd1000: data <= 8'h80;
            11'd1001: data <= 8'h80;
            11'd1002: data <= 8'h80;
            11'd1003: data <= 8'hBE;
            11'd1004: data <= 8'h80;
            11'd1005: data <= 8'hBE;
            11'd1006: data <= 8'h80;
            11'd1007: data <= 8'h80;
            11'd1008: data <= 8'h80;
            11'd1009: data <= 8'h90;
            11'd1010: data <= 8'h88;
            11'd1011: data <= 8'h84;
            11'd1012: data <= 8'h82;
            11'd1013: data <= 8'h84;
            11'd1014: data <= 8'h88;
            11'd1015: data <= 8'h90;
            11'd1016: data <= 8'h80;
            11'd1017: data <= 8'h9C;
            11'd1018: data <= 8'hA2;
            11'd1019: data <= 8'h84;
            11'd1020: data <= 8'h88;
            11'd1021: data <= 8'h88;
            11'd1022: data <= 8'h80;
            11'd1023: data <= 8'h88;
            11'd1024: data <= 8'h00;
            11'd1025: data <= 8'h1C;
            11'd1026: data <= 8'h22;
            11'd1027: data <= 8'h2A;
            11'd1028: data <= 8'h2E;
            11'd1029: data <= 8'h2C;
            11'd1030: data <= 8'h20;
            11'd1031: data <= 8'h1E;
            11'd1032: data <= 8'h00;
            11'd1033: data <= 8'h08;
            11'd1034: data <= 8'h14;
            11'd1035: data <= 8'h22;
            11'd1036: data <= 8'h22;
            11'd1037: data <= 8'h3E;
            11'd1038: data <= 8'h22;
            11'd1039: data <= 8'h22;
            11'd1040: data <= 8'h00;
            11'd1041: data <= 8'h3C;
            11'd1042: data <= 8'h22;
            11'd1043: data <= 8'h22;
            11'd1044: data <= 8'h3C;
            11'd1045: data <= 8'h22;
            11'd1046: data <= 8'h22;
            11'd1047: data <= 8'h3C;
            11'd1048: data <= 8'h00;
            11'd1049: data <= 8'h1C;
            11'd1050: data <= 8'h22;
            11'd1051: data <= 8'h20;
            11'd1052: data <= 8'h20;
            11'd1053: data <= 8'h20;
            11'd1054: data <= 8'h22;
            11'd1055: data <= 8'h1C;
            11'd1056: data <= 8'h00;
            11'd1057: data <= 8'h3C;
            11'd1058: data <= 8'h22;
            11'd1059: data <= 8'h22;
            11'd1060: data <= 8'h22;
            11'd1061: data <= 8'h22;
            11'd1062: data <= 8'h22;
            11'd1063: data <= 8'h3C;
            11'd1064: data <= 8'h00;
            11'd1065: data <= 8'h3E;
            11'd1066: data <= 8'h20;
            11'd1067: data <= 8'h20;
            11'd1068: data <= 8'h3C;
            11'd1069: data <= 8'h20;
            11'd1070: data <= 8'h20;
            11'd1071: data <= 8'h3E;
            11'd1072: data <= 8'h00;
            11'd1073: data <= 8'h3E;
            11'd1074: data <= 8'h20;
            11'd1075: data <= 8'h20;
            11'd1076: data <= 8'h3C;
            11'd1077: data <= 8'h20;
            11'd1078: data <= 8'h20;
            11'd1079: data <= 8'h20;
            11'd1080: data <= 8'h00;
            11'd1081: data <= 8'h1E;
            11'd1082: data <= 8'h20;
            11'd1083: data <= 8'h20;
            11'd1084: data <= 8'h20;
            11'd1085: data <= 8'h26;
            11'd1086: data <= 8'h22;
            11'd1087: data <= 8'h1E;
            11'd1088: data <= 8'h00;
            11'd1089: data <= 8'h22;
            11'd1090: data <= 8'h22;
            11'd1091: data <= 8'h22;
            11'd1092: data <= 8'h3E;
            11'd1093: data <= 8'h22;
            11'd1094: data <= 8'h22;
            11'd1095: data <= 8'h22;
            11'd1096: data <= 8'h00;
            11'd1097: data <= 8'h1C;
            11'd1098: data <= 8'h08;
            11'd1099: data <= 8'h08;
            11'd1100: data <= 8'h08;
            11'd1101: data <= 8'h08;
            11'd1102: data <= 8'h08;
            11'd1103: data <= 8'h1C;
            11'd1104: data <= 8'h00;
            11'd1105: data <= 8'h02;
            11'd1106: data <= 8'h02;
            11'd1107: data <= 8'h02;
            11'd1108: data <= 8'h02;
            11'd1109: data <= 8'h02;
            11'd1110: data <= 8'h22;
            11'd1111: data <= 8'h1C;
            11'd1112: data <= 8'h00;
            11'd1113: data <= 8'h22;
            11'd1114: data <= 8'h24;
            11'd1115: data <= 8'h28;
            11'd1116: data <= 8'h30;
            11'd1117: data <= 8'h28;
            11'd1118: data <= 8'h24;
            11'd1119: data <= 8'h22;
            11'd1120: data <= 8'h00;
            11'd1121: data <= 8'h20;
            11'd1122: data <= 8'h20;
            11'd1123: data <= 8'h20;
            11'd1124: data <= 8'h20;
            11'd1125: data <= 8'h20;
            11'd1126: data <= 8'h20;
            11'd1127: data <= 8'h3E;
            11'd1128: data <= 8'h00;
            11'd1129: data <= 8'h22;
            11'd1130: data <= 8'h36;
            11'd1131: data <= 8'h2A;
            11'd1132: data <= 8'h2A;
            11'd1133: data <= 8'h22;
            11'd1134: data <= 8'h22;
            11'd1135: data <= 8'h22;
            11'd1136: data <= 8'h00;
            11'd1137: data <= 8'h22;
            11'd1138: data <= 8'h22;
            11'd1139: data <= 8'h32;
            11'd1140: data <= 8'h2A;
            11'd1141: data <= 8'h26;
            11'd1142: data <= 8'h22;
            11'd1143: data <= 8'h22;
            11'd1144: data <= 8'h00;
            11'd1145: data <= 8'h1C;
            11'd1146: data <= 8'h22;
            11'd1147: data <= 8'h22;
            11'd1148: data <= 8'h22;
            11'd1149: data <= 8'h22;
            11'd1150: data <= 8'h22;
            11'd1151: data <= 8'h1C;
            11'd1152: data <= 8'h00;
            11'd1153: data <= 8'h3C;
            11'd1154: data <= 8'h22;
            11'd1155: data <= 8'h22;
            11'd1156: data <= 8'h3C;
            11'd1157: data <= 8'h20;
            11'd1158: data <= 8'h20;
            11'd1159: data <= 8'h20;
            11'd1160: data <= 8'h00;
            11'd1161: data <= 8'h1C;
            11'd1162: data <= 8'h22;
            11'd1163: data <= 8'h22;
            11'd1164: data <= 8'h22;
            11'd1165: data <= 8'h2A;
            11'd1166: data <= 8'h24;
            11'd1167: data <= 8'h1A;
            11'd1168: data <= 8'h00;
            11'd1169: data <= 8'h3C;
            11'd1170: data <= 8'h22;
            11'd1171: data <= 8'h22;
            11'd1172: data <= 8'h3C;
            11'd1173: data <= 8'h28;
            11'd1174: data <= 8'h24;
            11'd1175: data <= 8'h22;
            11'd1176: data <= 8'h00;
            11'd1177: data <= 8'h1C;
            11'd1178: data <= 8'h22;
            11'd1179: data <= 8'h20;
            11'd1180: data <= 8'h1C;
            11'd1181: data <= 8'h02;
            11'd1182: data <= 8'h22;
            11'd1183: data <= 8'h1C;
            11'd1184: data <= 8'h00;
            11'd1185: data <= 8'h3E;
            11'd1186: data <= 8'h08;
            11'd1187: data <= 8'h08;
            11'd1188: data <= 8'h08;
            11'd1189: data <= 8'h08;
            11'd1190: data <= 8'h08;
            11'd1191: data <= 8'h08;
            11'd1192: data <= 8'h00;
            11'd1193: data <= 8'h22;
            11'd1194: data <= 8'h22;
            11'd1195: data <= 8'h22;
            11'd1196: data <= 8'h22;
            11'd1197: data <= 8'h22;
            11'd1198: data <= 8'h22;
            11'd1199: data <= 8'h1C;
            11'd1200: data <= 8'h00;
            11'd1201: data <= 8'h22;
            11'd1202: data <= 8'h22;
            11'd1203: data <= 8'h22;
            11'd1204: data <= 8'h22;
            11'd1205: data <= 8'h22;
            11'd1206: data <= 8'h14;
            11'd1207: data <= 8'h08;
            11'd1208: data <= 8'h00;
            11'd1209: data <= 8'h22;
            11'd1210: data <= 8'h22;
            11'd1211: data <= 8'h22;
            11'd1212: data <= 8'h2A;
            11'd1213: data <= 8'h2A;
            11'd1214: data <= 8'h36;
            11'd1215: data <= 8'h22;
            11'd1216: data <= 8'h00;
            11'd1217: data <= 8'h22;
            11'd1218: data <= 8'h22;
            11'd1219: data <= 8'h14;
            11'd1220: data <= 8'h08;
            11'd1221: data <= 8'h14;
            11'd1222: data <= 8'h22;
            11'd1223: data <= 8'h22;
            11'd1224: data <= 8'h00;
            11'd1225: data <= 8'h22;
            11'd1226: data <= 8'h22;
            11'd1227: data <= 8'h14;
            11'd1228: data <= 8'h08;
            11'd1229: data <= 8'h08;
            11'd1230: data <= 8'h08;
            11'd1231: data <= 8'h08;
            11'd1232: data <= 8'h00;
            11'd1233: data <= 8'h3E;
            11'd1234: data <= 8'h02;
            11'd1235: data <= 8'h04;
            11'd1236: data <= 8'h08;
            11'd1237: data <= 8'h10;
            11'd1238: data <= 8'h20;
            11'd1239: data <= 8'h3E;
            11'd1240: data <= 8'h00;
            11'd1241: data <= 8'h3E;
            11'd1242: data <= 8'h30;
            11'd1243: data <= 8'h30;
            11'd1244: data <= 8'h30;
            11'd1245: data <= 8'h30;
            11'd1246: data <= 8'h30;
            11'd1247: data <= 8'h3E;
            11'd1248: data <= 8'h00;
            11'd1249: data <= 8'h00;
            11'd1250: data <= 8'h20;
            11'd1251: data <= 8'h10;
            11'd1252: data <= 8'h08;
            11'd1253: data <= 8'h04;
            11'd1254: data <= 8'h02;
            11'd1255: data <= 8'h00;
            11'd1256: data <= 8'h00;
            11'd1257: data <= 8'h3E;
            11'd1258: data <= 8'h06;
            11'd1259: data <= 8'h06;
            11'd1260: data <= 8'h06;
            11'd1261: data <= 8'h06;
            11'd1262: data <= 8'h06;
            11'd1263: data <= 8'h3E;
            11'd1264: data <= 8'h00;
            11'd1265: data <= 8'h00;
            11'd1266: data <= 8'h00;
            11'd1267: data <= 8'h08;
            11'd1268: data <= 8'h14;
            11'd1269: data <= 8'h22;
            11'd1270: data <= 8'h00;
            11'd1271: data <= 8'h00;
            11'd1272: data <= 8'h00;
            11'd1273: data <= 8'h00;
            11'd1274: data <= 8'h00;
            11'd1275: data <= 8'h00;
            11'd1276: data <= 8'h00;
            11'd1277: data <= 8'h00;
            11'd1278: data <= 8'h00;
            11'd1279: data <= 8'h3E;
            11'd1280: data <= 8'h00;
            11'd1281: data <= 8'h00;
            11'd1282: data <= 8'h00;
            11'd1283: data <= 8'h00;
            11'd1284: data <= 8'h00;
            11'd1285: data <= 8'h00;
            11'd1286: data <= 8'h00;
            11'd1287: data <= 8'h00;
            11'd1288: data <= 8'h00;
            11'd1289: data <= 8'h08;
            11'd1290: data <= 8'h08;
            11'd1291: data <= 8'h08;
            11'd1292: data <= 8'h08;
            11'd1293: data <= 8'h08;
            11'd1294: data <= 8'h00;
            11'd1295: data <= 8'h08;
            11'd1296: data <= 8'h00;
            11'd1297: data <= 8'h14;
            11'd1298: data <= 8'h14;
            11'd1299: data <= 8'h14;
            11'd1300: data <= 8'h00;
            11'd1301: data <= 8'h00;
            11'd1302: data <= 8'h00;
            11'd1303: data <= 8'h00;
            11'd1304: data <= 8'h00;
            11'd1305: data <= 8'h14;
            11'd1306: data <= 8'h14;
            11'd1307: data <= 8'h3E;
            11'd1308: data <= 8'h14;
            11'd1309: data <= 8'h3E;
            11'd1310: data <= 8'h14;
            11'd1311: data <= 8'h14;
            11'd1312: data <= 8'h00;
            11'd1313: data <= 8'h08;
            11'd1314: data <= 8'h1E;
            11'd1315: data <= 8'h28;
            11'd1316: data <= 8'h1C;
            11'd1317: data <= 8'h0A;
            11'd1318: data <= 8'h3C;
            11'd1319: data <= 8'h08;
            11'd1320: data <= 8'h00;
            11'd1321: data <= 8'h30;
            11'd1322: data <= 8'h32;
            11'd1323: data <= 8'h04;
            11'd1324: data <= 8'h08;
            11'd1325: data <= 8'h10;
            11'd1326: data <= 8'h26;
            11'd1327: data <= 8'h06;
            11'd1328: data <= 8'h00;
            11'd1329: data <= 8'h10;
            11'd1330: data <= 8'h28;
            11'd1331: data <= 8'h28;
            11'd1332: data <= 8'h10;
            11'd1333: data <= 8'h2A;
            11'd1334: data <= 8'h24;
            11'd1335: data <= 8'h1A;
            11'd1336: data <= 8'h00;
            11'd1337: data <= 8'h08;
            11'd1338: data <= 8'h08;
            11'd1339: data <= 8'h08;
            11'd1340: data <= 8'h00;
            11'd1341: data <= 8'h00;
            11'd1342: data <= 8'h00;
            11'd1343: data <= 8'h00;
            11'd1344: data <= 8'h00;
            11'd1345: data <= 8'h08;
            11'd1346: data <= 8'h10;
            11'd1347: data <= 8'h20;
            11'd1348: data <= 8'h20;
            11'd1349: data <= 8'h20;
            11'd1350: data <= 8'h10;
            11'd1351: data <= 8'h08;
            11'd1352: data <= 8'h00;
            11'd1353: data <= 8'h08;
            11'd1354: data <= 8'h04;
            11'd1355: data <= 8'h02;
            11'd1356: data <= 8'h02;
            11'd1357: data <= 8'h02;
            11'd1358: data <= 8'h04;
            11'd1359: data <= 8'h08;
            11'd1360: data <= 8'h00;
            11'd1361: data <= 8'h08;
            11'd1362: data <= 8'h2A;
            11'd1363: data <= 8'h1C;
            11'd1364: data <= 8'h08;
            11'd1365: data <= 8'h1C;
            11'd1366: data <= 8'h2A;
            11'd1367: data <= 8'h08;
            11'd1368: data <= 8'h00;
            11'd1369: data <= 8'h00;
            11'd1370: data <= 8'h08;
            11'd1371: data <= 8'h08;
            11'd1372: data <= 8'h3E;
            11'd1373: data <= 8'h08;
            11'd1374: data <= 8'h08;
            11'd1375: data <= 8'h00;
            11'd1376: data <= 8'h00;
            11'd1377: data <= 8'h00;
            11'd1378: data <= 8'h00;
            11'd1379: data <= 8'h00;
            11'd1380: data <= 8'h00;
            11'd1381: data <= 8'h08;
            11'd1382: data <= 8'h08;
            11'd1383: data <= 8'h10;
            11'd1384: data <= 8'h00;
            11'd1385: data <= 8'h00;
            11'd1386: data <= 8'h00;
            11'd1387: data <= 8'h00;
            11'd1388: data <= 8'h3E;
            11'd1389: data <= 8'h00;
            11'd1390: data <= 8'h00;
            11'd1391: data <= 8'h00;
            11'd1392: data <= 8'h00;
            11'd1393: data <= 8'h00;
            11'd1394: data <= 8'h00;
            11'd1395: data <= 8'h00;
            11'd1396: data <= 8'h00;
            11'd1397: data <= 8'h00;
            11'd1398: data <= 8'h00;
            11'd1399: data <= 8'h08;
            11'd1400: data <= 8'h00;
            11'd1401: data <= 8'h00;
            11'd1402: data <= 8'h02;
            11'd1403: data <= 8'h04;
            11'd1404: data <= 8'h08;
            11'd1405: data <= 8'h10;
            11'd1406: data <= 8'h20;
            11'd1407: data <= 8'h00;
            11'd1408: data <= 8'h00;
            11'd1409: data <= 8'h1C;
            11'd1410: data <= 8'h22;
            11'd1411: data <= 8'h26;
            11'd1412: data <= 8'h2A;
            11'd1413: data <= 8'h32;
            11'd1414: data <= 8'h22;
            11'd1415: data <= 8'h1C;
            11'd1416: data <= 8'h00;
            11'd1417: data <= 8'h08;
            11'd1418: data <= 8'h18;
            11'd1419: data <= 8'h08;
            11'd1420: data <= 8'h08;
            11'd1421: data <= 8'h08;
            11'd1422: data <= 8'h08;
            11'd1423: data <= 8'h1C;
            11'd1424: data <= 8'h00;
            11'd1425: data <= 8'h1C;
            11'd1426: data <= 8'h22;
            11'd1427: data <= 8'h02;
            11'd1428: data <= 8'h0C;
            11'd1429: data <= 8'h10;
            11'd1430: data <= 8'h20;
            11'd1431: data <= 8'h3E;
            11'd1432: data <= 8'h00;
            11'd1433: data <= 8'h3E;
            11'd1434: data <= 8'h02;
            11'd1435: data <= 8'h04;
            11'd1436: data <= 8'h0C;
            11'd1437: data <= 8'h02;
            11'd1438: data <= 8'h22;
            11'd1439: data <= 8'h1C;
            11'd1440: data <= 8'h00;
            11'd1441: data <= 8'h04;
            11'd1442: data <= 8'h0C;
            11'd1443: data <= 8'h14;
            11'd1444: data <= 8'h24;
            11'd1445: data <= 8'h3E;
            11'd1446: data <= 8'h04;
            11'd1447: data <= 8'h04;
            11'd1448: data <= 8'h00;
            11'd1449: data <= 8'h3E;
            11'd1450: data <= 8'h20;
            11'd1451: data <= 8'h3C;
            11'd1452: data <= 8'h02;
            11'd1453: data <= 8'h02;
            11'd1454: data <= 8'h22;
            11'd1455: data <= 8'h1C;
            11'd1456: data <= 8'h00;
            11'd1457: data <= 8'h0E;
            11'd1458: data <= 8'h10;
            11'd1459: data <= 8'h20;
            11'd1460: data <= 8'h3C;
            11'd1461: data <= 8'h22;
            11'd1462: data <= 8'h22;
            11'd1463: data <= 8'h1C;
            11'd1464: data <= 8'h00;
            11'd1465: data <= 8'h3E;
            11'd1466: data <= 8'h02;
            11'd1467: data <= 8'h04;
            11'd1468: data <= 8'h08;
            11'd1469: data <= 8'h10;
            11'd1470: data <= 8'h10;
            11'd1471: data <= 8'h10;
            11'd1472: data <= 8'h00;
            11'd1473: data <= 8'h1C;
            11'd1474: data <= 8'h22;
            11'd1475: data <= 8'h22;
            11'd1476: data <= 8'h1C;
            11'd1477: data <= 8'h22;
            11'd1478: data <= 8'h22;
            11'd1479: data <= 8'h1C;
            11'd1480: data <= 8'h00;
            11'd1481: data <= 8'h1C;
            11'd1482: data <= 8'h22;
            11'd1483: data <= 8'h22;
            11'd1484: data <= 8'h1E;
            11'd1485: data <= 8'h02;
            11'd1486: data <= 8'h04;
            11'd1487: data <= 8'h38;
            11'd1488: data <= 8'h00;
            11'd1489: data <= 8'h00;
            11'd1490: data <= 8'h00;
            11'd1491: data <= 8'h08;
            11'd1492: data <= 8'h00;
            11'd1493: data <= 8'h08;
            11'd1494: data <= 8'h00;
            11'd1495: data <= 8'h00;
            11'd1496: data <= 8'h00;
            11'd1497: data <= 8'h00;
            11'd1498: data <= 8'h00;
            11'd1499: data <= 8'h08;
            11'd1500: data <= 8'h00;
            11'd1501: data <= 8'h08;
            11'd1502: data <= 8'h08;
            11'd1503: data <= 8'h10;
            11'd1504: data <= 8'h00;
            11'd1505: data <= 8'h04;
            11'd1506: data <= 8'h08;
            11'd1507: data <= 8'h10;
            11'd1508: data <= 8'h20;
            11'd1509: data <= 8'h10;
            11'd1510: data <= 8'h08;
            11'd1511: data <= 8'h04;
            11'd1512: data <= 8'h00;
            11'd1513: data <= 8'h00;
            11'd1514: data <= 8'h00;
            11'd1515: data <= 8'h3E;
            11'd1516: data <= 8'h00;
            11'd1517: data <= 8'h3E;
            11'd1518: data <= 8'h00;
            11'd1519: data <= 8'h00;
            11'd1520: data <= 8'h00;
            11'd1521: data <= 8'h10;
            11'd1522: data <= 8'h08;
            11'd1523: data <= 8'h04;
            11'd1524: data <= 8'h02;
            11'd1525: data <= 8'h04;
            11'd1526: data <= 8'h08;
            11'd1527: data <= 8'h10;
            11'd1528: data <= 8'h00;
            11'd1529: data <= 8'h1C;
            11'd1530: data <= 8'h22;
            11'd1531: data <= 8'h04;
            11'd1532: data <= 8'h08;
            11'd1533: data <= 8'h08;
            11'd1534: data <= 8'h00;
            11'd1535: data <= 8'h08;
            11'd1536: data <= 8'h80;
            11'd1537: data <= 8'h9C;
            11'd1538: data <= 8'hA2;
            11'd1539: data <= 8'hAA;
            11'd1540: data <= 8'hAE;
            11'd1541: data <= 8'hAC;
            11'd1542: data <= 8'hA0;
            11'd1543: data <= 8'h9E;
            11'd1544: data <= 8'h80;
            11'd1545: data <= 8'h88;
            11'd1546: data <= 8'h94;
            11'd1547: data <= 8'hA2;
            11'd1548: data <= 8'hA2;
            11'd1549: data <= 8'hBE;
            11'd1550: data <= 8'hA2;
            11'd1551: data <= 8'hA2;
            11'd1552: data <= 8'h80;
            11'd1553: data <= 8'hBC;
            11'd1554: data <= 8'hA2;
            11'd1555: data <= 8'hA2;
            11'd1556: data <= 8'hBC;
            11'd1557: data <= 8'hA2;
            11'd1558: data <= 8'hA2;
            11'd1559: data <= 8'hBC;
            11'd1560: data <= 8'h80;
            11'd1561: data <= 8'h9C;
            11'd1562: data <= 8'hA2;
            11'd1563: data <= 8'hA0;
            11'd1564: data <= 8'hA0;
            11'd1565: data <= 8'hA0;
            11'd1566: data <= 8'hA2;
            11'd1567: data <= 8'h9C;
            11'd1568: data <= 8'h80;
            11'd1569: data <= 8'hBC;
            11'd1570: data <= 8'hA2;
            11'd1571: data <= 8'hA2;
            11'd1572: data <= 8'hA2;
            11'd1573: data <= 8'hA2;
            11'd1574: data <= 8'hA2;
            11'd1575: data <= 8'hBC;
            11'd1576: data <= 8'h80;
            11'd1577: data <= 8'hBE;
            11'd1578: data <= 8'hA0;
            11'd1579: data <= 8'hA0;
            11'd1580: data <= 8'hBC;
            11'd1581: data <= 8'hA0;
            11'd1582: data <= 8'hA0;
            11'd1583: data <= 8'hBE;
            11'd1584: data <= 8'h80;
            11'd1585: data <= 8'hBE;
            11'd1586: data <= 8'hA0;
            11'd1587: data <= 8'hA0;
            11'd1588: data <= 8'hBC;
            11'd1589: data <= 8'hA0;
            11'd1590: data <= 8'hA0;
            11'd1591: data <= 8'hA0;
            11'd1592: data <= 8'h80;
            11'd1593: data <= 8'h9E;
            11'd1594: data <= 8'hA0;
            11'd1595: data <= 8'hA0;
            11'd1596: data <= 8'hA0;
            11'd1597: data <= 8'hA6;
            11'd1598: data <= 8'hA2;
            11'd1599: data <= 8'h9E;
            11'd1600: data <= 8'h80;
            11'd1601: data <= 8'hA2;
            11'd1602: data <= 8'hA2;
            11'd1603: data <= 8'hA2;
            11'd1604: data <= 8'hBE;
            11'd1605: data <= 8'hA2;
            11'd1606: data <= 8'hA2;
            11'd1607: data <= 8'hA2;
            11'd1608: data <= 8'h80;
            11'd1609: data <= 8'h9C;
            11'd1610: data <= 8'h88;
            11'd1611: data <= 8'h88;
            11'd1612: data <= 8'h88;
            11'd1613: data <= 8'h88;
            11'd1614: data <= 8'h88;
            11'd1615: data <= 8'h9C;
            11'd1616: data <= 8'h80;
            11'd1617: data <= 8'h82;
            11'd1618: data <= 8'h82;
            11'd1619: data <= 8'h82;
            11'd1620: data <= 8'h82;
            11'd1621: data <= 8'h82;
            11'd1622: data <= 8'hA2;
            11'd1623: data <= 8'h9C;
            11'd1624: data <= 8'h80;
            11'd1625: data <= 8'hA2;
            11'd1626: data <= 8'hA4;
            11'd1627: data <= 8'hA8;
            11'd1628: data <= 8'hB0;
            11'd1629: data <= 8'hA8;
            11'd1630: data <= 8'hA4;
            11'd1631: data <= 8'hA2;
            11'd1632: data <= 8'h80;
            11'd1633: data <= 8'hA0;
            11'd1634: data <= 8'hA0;
            11'd1635: data <= 8'hA0;
            11'd1636: data <= 8'hA0;
            11'd1637: data <= 8'hA0;
            11'd1638: data <= 8'hA0;
            11'd1639: data <= 8'hBE;
            11'd1640: data <= 8'h80;
            11'd1641: data <= 8'hA2;
            11'd1642: data <= 8'hB6;
            11'd1643: data <= 8'hAA;
            11'd1644: data <= 8'hAA;
            11'd1645: data <= 8'hA2;
            11'd1646: data <= 8'hA2;
            11'd1647: data <= 8'hA2;
            11'd1648: data <= 8'h80;
            11'd1649: data <= 8'hA2;
            11'd1650: data <= 8'hA2;
            11'd1651: data <= 8'hB2;
            11'd1652: data <= 8'hAA;
            11'd1653: data <= 8'hA6;
            11'd1654: data <= 8'hA2;
            11'd1655: data <= 8'hA2;
            11'd1656: data <= 8'h80;
            11'd1657: data <= 8'h9C;
            11'd1658: data <= 8'hA2;
            11'd1659: data <= 8'hA2;
            11'd1660: data <= 8'hA2;
            11'd1661: data <= 8'hA2;
            11'd1662: data <= 8'hA2;
            11'd1663: data <= 8'h9C;
            11'd1664: data <= 8'h80;
            11'd1665: data <= 8'hBC;
            11'd1666: data <= 8'hA2;
            11'd1667: data <= 8'hA2;
            11'd1668: data <= 8'hBC;
            11'd1669: data <= 8'hA0;
            11'd1670: data <= 8'hA0;
            11'd1671: data <= 8'hA0;
            11'd1672: data <= 8'h80;
            11'd1673: data <= 8'h9C;
            11'd1674: data <= 8'hA2;
            11'd1675: data <= 8'hA2;
            11'd1676: data <= 8'hA2;
            11'd1677: data <= 8'hAA;
            11'd1678: data <= 8'hA4;
            11'd1679: data <= 8'h9A;
            11'd1680: data <= 8'h80;
            11'd1681: data <= 8'hBC;
            11'd1682: data <= 8'hA2;
            11'd1683: data <= 8'hA2;
            11'd1684: data <= 8'hBC;
            11'd1685: data <= 8'hA8;
            11'd1686: data <= 8'hA4;
            11'd1687: data <= 8'hA2;
            11'd1688: data <= 8'h80;
            11'd1689: data <= 8'h9C;
            11'd1690: data <= 8'hA2;
            11'd1691: data <= 8'hA0;
            11'd1692: data <= 8'h9C;
            11'd1693: data <= 8'h82;
            11'd1694: data <= 8'hA2;
            11'd1695: data <= 8'h9C;
            11'd1696: data <= 8'h80;
            11'd1697: data <= 8'hBE;
            11'd1698: data <= 8'h88;
            11'd1699: data <= 8'h88;
            11'd1700: data <= 8'h88;
            11'd1701: data <= 8'h88;
            11'd1702: data <= 8'h88;
            11'd1703: data <= 8'h88;
            11'd1704: data <= 8'h80;
            11'd1705: data <= 8'hA2;
            11'd1706: data <= 8'hA2;
            11'd1707: data <= 8'hA2;
            11'd1708: data <= 8'hA2;
            11'd1709: data <= 8'hA2;
            11'd1710: data <= 8'hA2;
            11'd1711: data <= 8'h9C;
            11'd1712: data <= 8'h80;
            11'd1713: data <= 8'hA2;
            11'd1714: data <= 8'hA2;
            11'd1715: data <= 8'hA2;
            11'd1716: data <= 8'hA2;
            11'd1717: data <= 8'hA2;
            11'd1718: data <= 8'h94;
            11'd1719: data <= 8'h88;
            11'd1720: data <= 8'h80;
            11'd1721: data <= 8'hA2;
            11'd1722: data <= 8'hA2;
            11'd1723: data <= 8'hA2;
            11'd1724: data <= 8'hAA;
            11'd1725: data <= 8'hAA;
            11'd1726: data <= 8'hB6;
            11'd1727: data <= 8'hA2;
            11'd1728: data <= 8'h80;
            11'd1729: data <= 8'hA2;
            11'd1730: data <= 8'hA2;
            11'd1731: data <= 8'h94;
            11'd1732: data <= 8'h88;
            11'd1733: data <= 8'h94;
            11'd1734: data <= 8'hA2;
            11'd1735: data <= 8'hA2;
            11'd1736: data <= 8'h80;
            11'd1737: data <= 8'hA2;
            11'd1738: data <= 8'hA2;
            11'd1739: data <= 8'h94;
            11'd1740: data <= 8'h88;
            11'd1741: data <= 8'h88;
            11'd1742: data <= 8'h88;
            11'd1743: data <= 8'h88;
            11'd1744: data <= 8'h80;
            11'd1745: data <= 8'hBE;
            11'd1746: data <= 8'h82;
            11'd1747: data <= 8'h84;
            11'd1748: data <= 8'h88;
            11'd1749: data <= 8'h90;
            11'd1750: data <= 8'hA0;
            11'd1751: data <= 8'hBE;
            11'd1752: data <= 8'h80;
            11'd1753: data <= 8'hBE;
            11'd1754: data <= 8'hB0;
            11'd1755: data <= 8'hB0;
            11'd1756: data <= 8'hB0;
            11'd1757: data <= 8'hB0;
            11'd1758: data <= 8'hB0;
            11'd1759: data <= 8'hBE;
            11'd1760: data <= 8'h80;
            11'd1761: data <= 8'h80;
            11'd1762: data <= 8'hA0;
            11'd1763: data <= 8'h90;
            11'd1764: data <= 8'h88;
            11'd1765: data <= 8'h84;
            11'd1766: data <= 8'h82;
            11'd1767: data <= 8'h80;
            11'd1768: data <= 8'h80;
            11'd1769: data <= 8'hBE;
            11'd1770: data <= 8'h86;
            11'd1771: data <= 8'h86;
            11'd1772: data <= 8'h86;
            11'd1773: data <= 8'h86;
            11'd1774: data <= 8'h86;
            11'd1775: data <= 8'hBE;
            11'd1776: data <= 8'h80;
            11'd1777: data <= 8'h80;
            11'd1778: data <= 8'h80;
            11'd1779: data <= 8'h88;
            11'd1780: data <= 8'h94;
            11'd1781: data <= 8'hA2;
            11'd1782: data <= 8'h80;
            11'd1783: data <= 8'h80;
            11'd1784: data <= 8'h80;
            11'd1785: data <= 8'h80;
            11'd1786: data <= 8'h80;
            11'd1787: data <= 8'h80;
            11'd1788: data <= 8'h80;
            11'd1789: data <= 8'h80;
            11'd1790: data <= 8'h80;
            11'd1791: data <= 8'hBE;
            11'd1792: data <= 8'h80;
            11'd1793: data <= 8'h80;
            11'd1794: data <= 8'h80;
            11'd1795: data <= 8'h80;
            11'd1796: data <= 8'h80;
            11'd1797: data <= 8'h80;
            11'd1798: data <= 8'h80;
            11'd1799: data <= 8'h80;
            11'd1800: data <= 8'h80;
            11'd1801: data <= 8'h88;
            11'd1802: data <= 8'h88;
            11'd1803: data <= 8'h88;
            11'd1804: data <= 8'h88;
            11'd1805: data <= 8'h88;
            11'd1806: data <= 8'h80;
            11'd1807: data <= 8'h88;
            11'd1808: data <= 8'h80;
            11'd1809: data <= 8'h94;
            11'd1810: data <= 8'h94;
            11'd1811: data <= 8'h94;
            11'd1812: data <= 8'h80;
            11'd1813: data <= 8'h80;
            11'd1814: data <= 8'h80;
            11'd1815: data <= 8'h80;
            11'd1816: data <= 8'h80;
            11'd1817: data <= 8'h94;
            11'd1818: data <= 8'h94;
            11'd1819: data <= 8'hBE;
            11'd1820: data <= 8'h94;
            11'd1821: data <= 8'hBE;
            11'd1822: data <= 8'h94;
            11'd1823: data <= 8'h94;
            11'd1824: data <= 8'h80;
            11'd1825: data <= 8'h88;
            11'd1826: data <= 8'h9E;
            11'd1827: data <= 8'hA8;
            11'd1828: data <= 8'h9C;
            11'd1829: data <= 8'h8A;
            11'd1830: data <= 8'hBC;
            11'd1831: data <= 8'h88;
            11'd1832: data <= 8'h80;
            11'd1833: data <= 8'hB0;
            11'd1834: data <= 8'hB2;
            11'd1835: data <= 8'h84;
            11'd1836: data <= 8'h88;
            11'd1837: data <= 8'h90;
            11'd1838: data <= 8'hA6;
            11'd1839: data <= 8'h86;
            11'd1840: data <= 8'h80;
            11'd1841: data <= 8'h90;
            11'd1842: data <= 8'hA8;
            11'd1843: data <= 8'hA8;
            11'd1844: data <= 8'h90;
            11'd1845: data <= 8'hAA;
            11'd1846: data <= 8'hA4;
            11'd1847: data <= 8'h9A;
            11'd1848: data <= 8'h80;
            11'd1849: data <= 8'h88;
            11'd1850: data <= 8'h88;
            11'd1851: data <= 8'h88;
            11'd1852: data <= 8'h80;
            11'd1853: data <= 8'h80;
            11'd1854: data <= 8'h80;
            11'd1855: data <= 8'h80;
            11'd1856: data <= 8'h80;
            11'd1857: data <= 8'h88;
            11'd1858: data <= 8'h90;
            11'd1859: data <= 8'hA0;
            11'd1860: data <= 8'hA0;
            11'd1861: data <= 8'hA0;
            11'd1862: data <= 8'h90;
            11'd1863: data <= 8'h88;
            11'd1864: data <= 8'h80;
            11'd1865: data <= 8'h88;
            11'd1866: data <= 8'h84;
            11'd1867: data <= 8'h82;
            11'd1868: data <= 8'h82;
            11'd1869: data <= 8'h82;
            11'd1870: data <= 8'h84;
            11'd1871: data <= 8'h88;
            11'd1872: data <= 8'h80;
            11'd1873: data <= 8'h88;
            11'd1874: data <= 8'hAA;
            11'd1875: data <= 8'h9C;
            11'd1876: data <= 8'h88;
            11'd1877: data <= 8'h9C;
            11'd1878: data <= 8'hAA;
            11'd1879: data <= 8'h88;
            11'd1880: data <= 8'h80;
            11'd1881: data <= 8'h80;
            11'd1882: data <= 8'h88;
            11'd1883: data <= 8'h88;
            11'd1884: data <= 8'hBE;
            11'd1885: data <= 8'h88;
            11'd1886: data <= 8'h88;
            11'd1887: data <= 8'h80;
            11'd1888: data <= 8'h80;
            11'd1889: data <= 8'h80;
            11'd1890: data <= 8'h80;
            11'd1891: data <= 8'h80;
            11'd1892: data <= 8'h80;
            11'd1893: data <= 8'h88;
            11'd1894: data <= 8'h88;
            11'd1895: data <= 8'h90;
            11'd1896: data <= 8'h80;
            11'd1897: data <= 8'h80;
            11'd1898: data <= 8'h80;
            11'd1899: data <= 8'h80;
            11'd1900: data <= 8'hBE;
            11'd1901: data <= 8'h80;
            11'd1902: data <= 8'h80;
            11'd1903: data <= 8'h80;
            11'd1904: data <= 8'h80;
            11'd1905: data <= 8'h80;
            11'd1906: data <= 8'h80;
            11'd1907: data <= 8'h80;
            11'd1908: data <= 8'h80;
            11'd1909: data <= 8'h80;
            11'd1910: data <= 8'h80;
            11'd1911: data <= 8'h88;
            11'd1912: data <= 8'h80;
            11'd1913: data <= 8'h80;
            11'd1914: data <= 8'h82;
            11'd1915: data <= 8'h84;
            11'd1916: data <= 8'h88;
            11'd1917: data <= 8'h90;
            11'd1918: data <= 8'hA0;
            11'd1919: data <= 8'h80;
            11'd1920: data <= 8'h80;
            11'd1921: data <= 8'h9C;
            11'd1922: data <= 8'hA2;
            11'd1923: data <= 8'hA6;
            11'd1924: data <= 8'hAA;
            11'd1925: data <= 8'hB2;
            11'd1926: data <= 8'hA2;
            11'd1927: data <= 8'h9C;
            11'd1928: data <= 8'h80;
            11'd1929: data <= 8'h88;
            11'd1930: data <= 8'h98;
            11'd1931: data <= 8'h88;
            11'd1932: data <= 8'h88;
            11'd1933: data <= 8'h88;
            11'd1934: data <= 8'h88;
            11'd1935: data <= 8'h9C;
            11'd1936: data <= 8'h80;
            11'd1937: data <= 8'h9C;
            11'd1938: data <= 8'hA2;
            11'd1939: data <= 8'h82;
            11'd1940: data <= 8'h8C;
            11'd1941: data <= 8'h90;
            11'd1942: data <= 8'hA0;
            11'd1943: data <= 8'hBE;
            11'd1944: data <= 8'h80;
            11'd1945: data <= 8'hBE;
            11'd1946: data <= 8'h82;
            11'd1947: data <= 8'h84;
            11'd1948: data <= 8'h8C;
            11'd1949: data <= 8'h82;
            11'd1950: data <= 8'hA2;
            11'd1951: data <= 8'h9C;
            11'd1952: data <= 8'h80;
            11'd1953: data <= 8'h84;
            11'd1954: data <= 8'h8C;
            11'd1955: data <= 8'h94;
            11'd1956: data <= 8'hA4;
            11'd1957: data <= 8'hBE;
            11'd1958: data <= 8'h84;
            11'd1959: data <= 8'h84;
            11'd1960: data <= 8'h80;
            11'd1961: data <= 8'hBE;
            11'd1962: data <= 8'hA0;
            11'd1963: data <= 8'hBC;
            11'd1964: data <= 8'h82;
            11'd1965: data <= 8'h82;
            11'd1966: data <= 8'hA2;
            11'd1967: data <= 8'h9C;
            11'd1968: data <= 8'h80;
            11'd1969: data <= 8'h8E;
            11'd1970: data <= 8'h90;
            11'd1971: data <= 8'hA0;
            11'd1972: data <= 8'hBC;
            11'd1973: data <= 8'hA2;
            11'd1974: data <= 8'hA2;
            11'd1975: data <= 8'h9C;
            11'd1976: data <= 8'h80;
            11'd1977: data <= 8'hBE;
            11'd1978: data <= 8'h82;
            11'd1979: data <= 8'h84;
            11'd1980: data <= 8'h88;
            11'd1981: data <= 8'h90;
            11'd1982: data <= 8'h90;
            11'd1983: data <= 8'h90;
            11'd1984: data <= 8'h80;
            11'd1985: data <= 8'h9C;
            11'd1986: data <= 8'hA2;
            11'd1987: data <= 8'hA2;
            11'd1988: data <= 8'h9C;
            11'd1989: data <= 8'hA2;
            11'd1990: data <= 8'hA2;
            11'd1991: data <= 8'h9C;
            11'd1992: data <= 8'h80;
            11'd1993: data <= 8'h9C;
            11'd1994: data <= 8'hA2;
            11'd1995: data <= 8'hA2;
            11'd1996: data <= 8'h9E;
            11'd1997: data <= 8'h82;
            11'd1998: data <= 8'h84;
            11'd1999: data <= 8'hB8;
            11'd2000: data <= 8'h80;
            11'd2001: data <= 8'h80;
            11'd2002: data <= 8'h80;
            11'd2003: data <= 8'h88;
            11'd2004: data <= 8'h80;
            11'd2005: data <= 8'h88;
            11'd2006: data <= 8'h80;
            11'd2007: data <= 8'h80;
            11'd2008: data <= 8'h80;
            11'd2009: data <= 8'h80;
            11'd2010: data <= 8'h80;
            11'd2011: data <= 8'h88;
            11'd2012: data <= 8'h80;
            11'd2013: data <= 8'h88;
            11'd2014: data <= 8'h88;
            11'd2015: data <= 8'h90;
            11'd2016: data <= 8'h80;
            11'd2017: data <= 8'h84;
            11'd2018: data <= 8'h88;
            11'd2019: data <= 8'h90;
            11'd2020: data <= 8'hA0;
            11'd2021: data <= 8'h90;
            11'd2022: data <= 8'h88;
            11'd2023: data <= 8'h84;
            11'd2024: data <= 8'h80;
            11'd2025: data <= 8'h80;
            11'd2026: data <= 8'h80;
            11'd2027: data <= 8'hBE;
            11'd2028: data <= 8'h80;
            11'd2029: data <= 8'hBE;
            11'd2030: data <= 8'h80;
            11'd2031: data <= 8'h80;
            11'd2032: data <= 8'h80;
            11'd2033: data <= 8'h90;
            11'd2034: data <= 8'h88;
            11'd2035: data <= 8'h84;
            11'd2036: data <= 8'h82;
            11'd2037: data <= 8'h84;
            11'd2038: data <= 8'h88;
            11'd2039: data <= 8'h90;
            11'd2040: data <= 8'h80;
            11'd2041: data <= 8'h9C;
            11'd2042: data <= 8'hA2;
            11'd2043: data <= 8'h84;
            11'd2044: data <= 8'h88;
            11'd2045: data <= 8'h88;
            11'd2046: data <= 8'h80;
            11'd2047: data <= 8'h88;
            default: data <= 8'h00;
        endcase
    end
endmodule
