`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/17/2025 08:23:27 PM
// Design Name: 
// Module Name: rom
// Project Name: 
// Target Devices: 
//////////////////////////////////////////////////////////////////////////////////



////-------------------------------------------------------------------------------------------------
module monitor_rom
//-------------------------------------------------------------------------------------------------
#
(
	parameter DW = 8,
	parameter AW = 14
)
(
	input  wire         clock,
	input  wire         ce,
	output reg [DW-1:0] data_out,
	input  wire[AW-1:0] a
);
//-------------------------------------------------------------------------------------------------

reg[DW-1:0] d[(2**AW)-1:0];
initial $readmemb("Apple II ROM Pages F8-FF - 341-0004 - Original Monitor.bin", d);

always @(posedge clock) if(ce) data_out<= d[a];

//-------------------------------------------------------------------------------------------------
endmodule
////-------------------------------------------------------------------------------------------------
